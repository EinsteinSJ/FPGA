-- PLL_3orden_change_GN_PLL_3orden_change_PLL_ab_dq.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PLL_3orden_change_GN_PLL_3orden_change_PLL_ab_dq is
	port (
		a       : in  std_logic_vector(13 downto 0) := (others => '0'); --       a.wire
		alpha_o : in  std_logic_vector(9 downto 0)  := (others => '0'); -- alpha_o.wire
		b       : in  std_logic_vector(13 downto 0) := (others => '0'); --       b.wire
		Vd      : out std_logic_vector(13 downto 0);                    --      Vd.wire
		Clock   : in  std_logic                     := '0';             --   Clock.clk
		aclr    : in  std_logic                     := '0';             --        .reset
		Vq      : out std_logic_vector(13 downto 0)                     --      Vq.wire
	);
end entity PLL_3orden_change_GN_PLL_3orden_change_PLL_ab_dq;

architecture rtl of PLL_3orden_change_GN_PLL_3orden_change_PLL_ab_dq is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_multiplier_GNXOJHAPZV is
		generic (
			aWidth                         : natural := 8;
			Signed                         : natural := 0;
			bWidth                         : natural := 8;
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			pipeline                       : integer := 0;
			OutputLsb                      : integer := 0;
			OutputMsb                      : integer := 8
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GNXOJHAPZV;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_port_GNBOOX3JQY is
		port (
			input  : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNBOOX3JQY;

	component alt_dspbuilder_pipelined_adder_GN4HTUTWRG is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GN4HTUTWRG;

	component alt_dspbuilder_pipelined_adder_GNY2JEH574 is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNY2JEH574;

	component alt_dspbuilder_port_GNSSYS4J5R is
		port (
			input  : in  std_logic_vector(9 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(9 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNSSYS4J5R;

	component PLL_3orden_change_GN_PLL_3orden_change_PLL_ab_dq_SIN_COS is
		port (
			alpha_o : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- wire
			Clock   : in  std_logic                     := 'X';             -- clk
			aclr    : in  std_logic                     := 'X';             -- reset
			SIN1    : out std_logic_vector(13 downto 0);                    -- wire
			COS1    : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component PLL_3orden_change_GN_PLL_3orden_change_PLL_ab_dq_SIN_COS;

	signal multiplier2user_aclrgnd_output_wire             : std_logic;                     -- Multiplier2user_aclrGND:output -> Multiplier2:user_aclr
	signal multiplier2enavcc_output_wire                   : std_logic;                     -- Multiplier2enaVCC:output -> Multiplier2:ena
	signal multiplier1user_aclrgnd_output_wire             : std_logic;                     -- Multiplier1user_aclrGND:output -> Multiplier1:user_aclr
	signal multiplier1enavcc_output_wire                   : std_logic;                     -- Multiplier1enaVCC:output -> Multiplier1:ena
	signal multiplier3user_aclrgnd_output_wire             : std_logic;                     -- Multiplier3user_aclrGND:output -> Multiplier3:user_aclr
	signal multiplier3enavcc_output_wire                   : std_logic;                     -- Multiplier3enaVCC:output -> Multiplier3:ena
	signal multiplieruser_aclrgnd_output_wire              : std_logic;                     -- Multiplieruser_aclrGND:output -> Multiplier:user_aclr
	signal multiplierenavcc_output_wire                    : std_logic;                     -- MultiplierenaVCC:output -> Multiplier:ena
	signal pipelined_adderuser_aclrgnd_output_wire         : std_logic;                     -- Pipelined_Adderuser_aclrGND:output -> Pipelined_Adder:user_aclr
	signal pipelined_adderenavcc_output_wire               : std_logic;                     -- Pipelined_AdderenaVCC:output -> Pipelined_Adder:ena
	signal pipelined_adder1user_aclrgnd_output_wire        : std_logic;                     -- Pipelined_Adder1user_aclrGND:output -> Pipelined_Adder1:user_aclr
	signal pipelined_adder1enavcc_output_wire              : std_logic;                     -- Pipelined_Adder1enaVCC:output -> Pipelined_Adder1:ena
	signal a_0_output_wire                                 : std_logic_vector(13 downto 0); -- a_0:output -> [Multiplier3:dataa, Multiplier:dataa]
	signal b_0_output_wire                                 : std_logic_vector(13 downto 0); -- b_0:output -> [Multiplier1:dataa, Multiplier2:dataa]
	signal multiplier_result_wire                          : std_logic_vector(13 downto 0); -- Multiplier:result -> Pipelined_Adder:dataa
	signal multiplier1_result_wire                         : std_logic_vector(13 downto 0); -- Multiplier1:result -> Pipelined_Adder:datab
	signal multiplier2_result_wire                         : std_logic_vector(13 downto 0); -- Multiplier2:result -> Pipelined_Adder1:dataa
	signal multiplier3_result_wire                         : std_logic_vector(13 downto 0); -- Multiplier3:result -> Pipelined_Adder1:datab
	signal alpha_o_0_output_wire                           : std_logic_vector(9 downto 0);  -- alpha_o_0:output -> PLL_3orden_change_PLL_ab_dq_SIN_COS_0:alpha_o
	signal pll_3orden_change_pll_ab_dq_sin_cos_0_sin1_wire : std_logic_vector(13 downto 0); -- PLL_3orden_change_PLL_ab_dq_SIN_COS_0:SIN1 -> [Multiplier1:datab, Multiplier3:datab]
	signal pll_3orden_change_pll_ab_dq_sin_cos_0_cos1_wire : std_logic_vector(13 downto 0); -- PLL_3orden_change_PLL_ab_dq_SIN_COS_0:COS1 -> [Multiplier2:datab, Multiplier:datab]
	signal pipelined_adder_result_wire                     : std_logic_vector(13 downto 0); -- Pipelined_Adder:result -> Vd_0:input
	signal pipelined_adder1_result_wire                    : std_logic_vector(13 downto 0); -- Pipelined_Adder1:result -> Vq_0:input
	signal clock_0_clock_output_clk                        : std_logic;                     -- Clock_0:clock_out -> [Multiplier1:clock, Multiplier2:clock, Multiplier3:clock, Multiplier:clock, PLL_3orden_change_PLL_ab_dq_SIN_COS_0:Clock, Pipelined_Adder1:clock, Pipelined_Adder:clock]
	signal clock_0_clock_output_reset                      : std_logic;                     -- Clock_0:aclr_out -> [Multiplier1:aclr, Multiplier2:aclr, Multiplier3:aclr, Multiplier:aclr, PLL_3orden_change_PLL_ab_dq_SIN_COS_0:aclr, Pipelined_Adder1:aclr, Pipelined_Adder:aclr]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	multiplier2 : component alt_dspbuilder_multiplier_GNXOJHAPZV
		generic map (
			aWidth                         => 14,
			Signed                         => 1,
			bWidth                         => 14,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 1,
			OutputLsb                      => 12,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,                        -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                      --           .reset
			dataa     => b_0_output_wire,                                 --      dataa.wire
			datab     => pll_3orden_change_pll_ab_dq_sin_cos_0_cos1_wire, --      datab.wire
			result    => multiplier2_result_wire,                         --     result.wire
			user_aclr => multiplier2user_aclrgnd_output_wire,             --  user_aclr.wire
			ena       => multiplier2enavcc_output_wire                    --        ena.wire
		);

	multiplier2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier2user_aclrgnd_output_wire  -- output.wire
		);

	multiplier2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplier2enavcc_output_wire  -- output.wire
		);

	a_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => a,               --  input.wire
			output => a_0_output_wire  -- output.wire
		);

	multiplier1 : component alt_dspbuilder_multiplier_GNXOJHAPZV
		generic map (
			aWidth                         => 14,
			Signed                         => 1,
			bWidth                         => 14,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 1,
			OutputLsb                      => 12,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,                        -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                      --           .reset
			dataa     => b_0_output_wire,                                 --      dataa.wire
			datab     => pll_3orden_change_pll_ab_dq_sin_cos_0_sin1_wire, --      datab.wire
			result    => multiplier1_result_wire,                         --     result.wire
			user_aclr => multiplier1user_aclrgnd_output_wire,             --  user_aclr.wire
			ena       => multiplier1enavcc_output_wire                    --        ena.wire
		);

	multiplier1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier1user_aclrgnd_output_wire  -- output.wire
		);

	multiplier1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplier1enavcc_output_wire  -- output.wire
		);

	b_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => b,               --  input.wire
			output => b_0_output_wire  -- output.wire
		);

	multiplier3 : component alt_dspbuilder_multiplier_GNXOJHAPZV
		generic map (
			aWidth                         => 14,
			Signed                         => 1,
			bWidth                         => 14,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 1,
			OutputLsb                      => 12,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,                        -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                      --           .reset
			dataa     => a_0_output_wire,                                 --      dataa.wire
			datab     => pll_3orden_change_pll_ab_dq_sin_cos_0_sin1_wire, --      datab.wire
			result    => multiplier3_result_wire,                         --     result.wire
			user_aclr => multiplier3user_aclrgnd_output_wire,             --  user_aclr.wire
			ena       => multiplier3enavcc_output_wire                    --        ena.wire
		);

	multiplier3user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier3user_aclrgnd_output_wire  -- output.wire
		);

	multiplier3enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplier3enavcc_output_wire  -- output.wire
		);

	multiplier : component alt_dspbuilder_multiplier_GNXOJHAPZV
		generic map (
			aWidth                         => 14,
			Signed                         => 1,
			bWidth                         => 14,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 1,
			OutputLsb                      => 12,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,                        -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                      --           .reset
			dataa     => a_0_output_wire,                                 --      dataa.wire
			datab     => pll_3orden_change_pll_ab_dq_sin_cos_0_cos1_wire, --      datab.wire
			result    => multiplier_result_wire,                          --     result.wire
			user_aclr => multiplieruser_aclrgnd_output_wire,              --  user_aclr.wire
			ena       => multiplierenavcc_output_wire                     --        ena.wire
		);

	multiplieruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplieruser_aclrgnd_output_wire  -- output.wire
		);

	multiplierenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplierenavcc_output_wire  -- output.wire
		);

	pipelined_adder : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 14
		)
		port map (
			clock     => clock_0_clock_output_clk,                -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,              --           .reset
			dataa     => multiplier_result_wire,                  --      dataa.wire
			datab     => multiplier1_result_wire,                 --      datab.wire
			result    => pipelined_adder_result_wire,             --     result.wire
			user_aclr => pipelined_adderuser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adderenavcc_output_wire        --        ena.wire
		);

	pipelined_adderuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adderuser_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adderenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adderenavcc_output_wire  -- output.wire
		);

	pipelined_adder1 : component alt_dspbuilder_pipelined_adder_GNY2JEH574
		generic map (
			pipeline => 0,
			width    => 14
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => multiplier2_result_wire,                  --      dataa.wire
			datab     => multiplier3_result_wire,                  --      datab.wire
			result    => pipelined_adder1_result_wire,             --     result.wire
			user_aclr => pipelined_adder1user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder1enavcc_output_wire        --        ena.wire
		);

	pipelined_adder1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder1user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder1enavcc_output_wire  -- output.wire
		);

	vq_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => pipelined_adder1_result_wire, --  input.wire
			output => Vq                            -- output.wire
		);

	alpha_o_0 : component alt_dspbuilder_port_GNSSYS4J5R
		port map (
			input  => alpha_o,               --  input.wire
			output => alpha_o_0_output_wire  -- output.wire
		);

	pll_3orden_change_pll_ab_dq_sin_cos_0 : component PLL_3orden_change_GN_PLL_3orden_change_PLL_ab_dq_SIN_COS
		port map (
			alpha_o => alpha_o_0_output_wire,                           -- alpha_o.wire
			Clock   => clock_0_clock_output_clk,                        --   Clock.clk
			aclr    => clock_0_clock_output_reset,                      --        .reset
			SIN1    => pll_3orden_change_pll_ab_dq_sin_cos_0_sin1_wire, --    SIN1.wire
			COS1    => pll_3orden_change_pll_ab_dq_sin_cos_0_cos1_wire  --    COS1.wire
		);

	vd_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => pipelined_adder_result_wire, --  input.wire
			output => Vd                           -- output.wire
		);

end architecture rtl; -- of PLL_3orden_change_GN_PLL_3orden_change_PLL_ab_dq
