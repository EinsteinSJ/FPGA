-- PLL_3orden_change_GN_PLL_3orden_change_PLL_PI_z.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PLL_3orden_change_GN_PLL_3orden_change_PLL_PI_z is
	port (
		Clock     : in  std_logic                     := '0';             --     Clock.clk
		aclr      : in  std_logic                     := '0';             --          .reset
		Vd        : in  std_logic_vector(13 downto 0) := (others => '0'); --        Vd.wire
		Wo_ref    : in  std_logic_vector(13 downto 0) := (others => '0'); --    Wo_ref.wire
		wo        : out std_logic_vector(17 downto 0);                    --        wo.wire
		Ts        : in  std_logic_vector(31 downto 0) := (others => '0'); --        Ts.wire
		CLK_60KHz : in  std_logic                     := '0'              -- CLK_60KHz.wire
	);
end entity PLL_3orden_change_GN_PLL_3orden_change_PLL_PI_z;

architecture rtl of PLL_3orden_change_GN_PLL_3orden_change_PLL_PI_z is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_cast_GNF7MCRHPM is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNF7MCRHPM;

	component alt_dspbuilder_cast_GND47QX5DY is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GND47QX5DY;

	component alt_dspbuilder_multiplier_GNWKYNVRFY is
		generic (
			aWidth                         : natural := 8;
			Signed                         : natural := 0;
			bWidth                         : natural := 8;
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			pipeline                       : integer := 0;
			OutputLsb                      : integer := 0;
			OutputMsb                      : integer := 8
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GNWKYNVRFY;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_constant_GN6EHA4QWH is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(17 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GN6EHA4QWH;

	component alt_dspbuilder_pipelined_adder_GN4HTUTWRG is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GN4HTUTWRG;

	component PLL_3orden_change_GN_PLL_3orden_change_PLL_PI_z_1_sv2 is
		port (
			Clock   : in  std_logic                     := 'X';             -- clk
			aclr    : in  std_logic                     := 'X';             -- reset
			CLK_60K : in  std_logic                     := 'X';             -- wire
			Ts      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			Vd      : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			E       : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component PLL_3orden_change_GN_PLL_3orden_change_PLL_PI_z_1_sv2;

	component alt_dspbuilder_port_GNBOOX3JQY is
		port (
			input  : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNBOOX3JQY;

	component alt_dspbuilder_port_GN2CABCRLL is
		port (
			input  : in  std_logic_vector(17 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(17 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GN2CABCRLL;

	component alt_dspbuilder_cast_GNBBMDRQ7A is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNBBMDRQ7A;

	component alt_dspbuilder_cast_GN6DTGWIDG is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(17 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(17 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN6DTGWIDG;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component alt_dspbuilder_cast_GNLZYLEWIQ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(17 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(17 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNLZYLEWIQ;

	component alt_dspbuilder_cast_GNSPENWJQH is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNSPENWJQH;

	component alt_dspbuilder_cast_GNQP67JAWW is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNQP67JAWW;

	component alt_dspbuilder_cast_GNXY6JKR5E is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNXY6JKR5E;

	component alt_dspbuilder_cast_GNRB4ECDTY is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(17 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNRB4ECDTY;

	component alt_dspbuilder_cast_GNCDTXOZMF is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(17 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNCDTXOZMF;

	component alt_dspbuilder_cast_GNWHGOINAS is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNWHGOINAS;

	signal multiplier1user_aclrgnd_output_wire       : std_logic;                     -- Multiplier1user_aclrGND:output -> Multiplier1:user_aclr
	signal multiplier1enavcc_output_wire             : std_logic;                     -- Multiplier1enaVCC:output -> Multiplier1:ena
	signal pipelined_adderuser_aclrgnd_output_wire   : std_logic;                     -- Pipelined_Adderuser_aclrGND:output -> Pipelined_Adder:user_aclr
	signal pipelined_adderenavcc_output_wire         : std_logic;                     -- Pipelined_AdderenaVCC:output -> Pipelined_Adder:ena
	signal pipelined_adder1user_aclrgnd_output_wire  : std_logic;                     -- Pipelined_Adder1user_aclrGND:output -> Pipelined_Adder1:user_aclr
	signal pipelined_adder1enavcc_output_wire        : std_logic;                     -- Pipelined_Adder1enaVCC:output -> Pipelined_Adder1:ena
	signal vd_0_output_wire                          : std_logic_vector(13 downto 0); -- Vd_0:output -> [PLL_3orden_change_PLL_PI_z_1_sv2_0:Vd, cast7:input]
	signal clk_60khz_0_output_wire                   : std_logic;                     -- CLK_60KHz_0:output -> PLL_3orden_change_PLL_PI_z_1_sv2_0:CLK_60K
	signal ts_0_output_wire                          : std_logic_vector(31 downto 0); -- Ts_0:output -> PLL_3orden_change_PLL_PI_z_1_sv2_0:Ts
	signal bus_conversion5_output_wire               : std_logic_vector(17 downto 0); -- Bus_Conversion5:output -> Multiplier1:dataa
	signal k2_output_wire                            : std_logic_vector(17 downto 0); -- K2:output -> Multiplier1:datab
	signal multiplier1_result_wire                   : std_logic_vector(31 downto 0); -- Multiplier1:result -> Bus_Conversion6:input
	signal bus_conversion2_output_wire               : std_logic_vector(31 downto 0); -- Bus_Conversion2:output -> Pipelined_Adder:dataa
	signal bus_conversion3_output_wire               : std_logic_vector(31 downto 0); -- Bus_Conversion3:output -> Pipelined_Adder:datab
	signal bus_conversion4_output_wire               : std_logic_vector(31 downto 0); -- Bus_Conversion4:output -> Pipelined_Adder1:dataa
	signal bus_conversion6_output_wire               : std_logic_vector(31 downto 0); -- Bus_Conversion6:output -> Pipelined_Adder1:datab
	signal bus_conversion1_output_wire               : std_logic_vector(31 downto 0); -- Bus_Conversion1:output -> x0_5:input
	signal bus_conversion7_output_wire               : std_logic_vector(17 downto 0); -- Bus_Conversion7:output -> wo_0:input
	signal cast7_output_wire                         : std_logic_vector(31 downto 0); -- cast7:output -> Bus_Conversion1:input
	signal pll_3orden_change_pll_pi_z_1_sv2_0_e_wire : std_logic_vector(31 downto 0); -- PLL_3orden_change_PLL_PI_z_1_sv2_0:E -> cast8:input
	signal cast8_output_wire                         : std_logic_vector(31 downto 0); -- cast8:output -> Bus_Conversion2:input
	signal wo_ref_0_output_wire                      : std_logic_vector(13 downto 0); -- Wo_ref_0:output -> cast9:input
	signal cast9_output_wire                         : std_logic_vector(31 downto 0); -- cast9:output -> Bus_Conversion4:input
	signal pipelined_adder_result_wire               : std_logic_vector(31 downto 0); -- Pipelined_Adder:result -> cast10:input
	signal cast10_output_wire                        : std_logic_vector(17 downto 0); -- cast10:output -> Bus_Conversion5:input
	signal pipelined_adder1_result_wire              : std_logic_vector(31 downto 0); -- Pipelined_Adder1:result -> cast11:input
	signal cast11_output_wire                        : std_logic_vector(17 downto 0); -- cast11:output -> Bus_Conversion7:input
	signal x0_5_output_wire                          : std_logic_vector(31 downto 0); -- x0_5:output -> cast12:input
	signal cast12_output_wire                        : std_logic_vector(31 downto 0); -- cast12:output -> Bus_Conversion3:input
	signal clock_0_clock_output_clk                  : std_logic;                     -- Clock_0:clock_out -> [Multiplier1:clock, PLL_3orden_change_PLL_PI_z_1_sv2_0:Clock, Pipelined_Adder1:clock, Pipelined_Adder:clock]
	signal clock_0_clock_output_reset                : std_logic;                     -- Clock_0:aclr_out -> [Multiplier1:aclr, PLL_3orden_change_PLL_PI_z_1_sv2_0:aclr, Pipelined_Adder1:aclr, Pipelined_Adder:aclr]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	bus_conversion4 : component alt_dspbuilder_cast_GNF7MCRHPM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast9_output_wire,           --  input.wire
			output => bus_conversion4_output_wire  -- output.wire
		);

	bus_conversion3 : component alt_dspbuilder_cast_GND47QX5DY
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast12_output_wire,          --  input.wire
			output => bus_conversion3_output_wire  -- output.wire
		);

	multiplier1 : component alt_dspbuilder_multiplier_GNWKYNVRFY
		generic map (
			aWidth                         => 18,
			Signed                         => 1,
			bWidth                         => 18,
			DEDICATED_MULTIPLIER_CIRCUITRY => "YES",
			pipeline                       => 1,
			OutputLsb                      => 3,
			OutputMsb                      => 34
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			dataa     => bus_conversion5_output_wire,         --      dataa.wire
			datab     => k2_output_wire,                      --      datab.wire
			result    => multiplier1_result_wire,             --     result.wire
			user_aclr => multiplier1user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => multiplier1enavcc_output_wire        --        ena.wire
		);

	multiplier1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier1user_aclrgnd_output_wire  -- output.wire
		);

	multiplier1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplier1enavcc_output_wire  -- output.wire
		);

	bus_conversion2 : component alt_dspbuilder_cast_GND47QX5DY
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast8_output_wire,           --  input.wire
			output => bus_conversion2_output_wire  -- output.wire
		);

	bus_conversion1 : component alt_dspbuilder_cast_GND47QX5DY
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast7_output_wire,           --  input.wire
			output => bus_conversion1_output_wire  -- output.wire
		);

	clk_60khz_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => CLK_60KHz,               --  input.wire
			output => clk_60khz_0_output_wire  -- output.wire
		);

	k2 : component alt_dspbuilder_constant_GN6EHA4QWH
		generic map (
			BitPattern => "010001101010111000",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 18
		)
		port map (
			output => k2_output_wire  -- output.wire
		);

	pipelined_adder : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 32
		)
		port map (
			clock     => clock_0_clock_output_clk,                -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,              --           .reset
			dataa     => bus_conversion2_output_wire,             --      dataa.wire
			datab     => bus_conversion3_output_wire,             --      datab.wire
			result    => pipelined_adder_result_wire,             --     result.wire
			user_aclr => pipelined_adderuser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adderenavcc_output_wire        --        ena.wire
		);

	pipelined_adderuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adderuser_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adderenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adderenavcc_output_wire  -- output.wire
		);

	pll_3orden_change_pll_pi_z_1_sv2_0 : component PLL_3orden_change_GN_PLL_3orden_change_PLL_PI_z_1_sv2
		port map (
			Clock   => clock_0_clock_output_clk,                  --   Clock.clk
			aclr    => clock_0_clock_output_reset,                --        .reset
			CLK_60K => clk_60khz_0_output_wire,                   -- CLK_60K.wire
			Ts      => ts_0_output_wire,                          --      Ts.wire
			Vd      => vd_0_output_wire,                          --      Vd.wire
			E       => pll_3orden_change_pll_pi_z_1_sv2_0_e_wire  --       E.wire
		);

	vd_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => Vd,               --  input.wire
			output => vd_0_output_wire  -- output.wire
		);

	wo_ref_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => Wo_ref,               --  input.wire
			output => wo_ref_0_output_wire  -- output.wire
		);

	wo_0 : component alt_dspbuilder_port_GN2CABCRLL
		port map (
			input  => bus_conversion7_output_wire, --  input.wire
			output => wo                           -- output.wire
		);

	x0_5 : component alt_dspbuilder_cast_GNBBMDRQ7A
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => bus_conversion1_output_wire, --  input.wire
			output => x0_5_output_wire             -- output.wire
		);

	pipelined_adder1 : component alt_dspbuilder_pipelined_adder_GN4HTUTWRG
		generic map (
			pipeline => 0,
			width    => 32
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => bus_conversion4_output_wire,              --      dataa.wire
			datab     => bus_conversion6_output_wire,              --      datab.wire
			result    => pipelined_adder1_result_wire,             --     result.wire
			user_aclr => pipelined_adder1user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder1enavcc_output_wire        --        ena.wire
		);

	pipelined_adder1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder1user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder1enavcc_output_wire  -- output.wire
		);

	bus_conversion7 : component alt_dspbuilder_cast_GN6DTGWIDG
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast11_output_wire,          --  input.wire
			output => bus_conversion7_output_wire  -- output.wire
		);

	bus_conversion6 : component alt_dspbuilder_cast_GNF7MCRHPM
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier1_result_wire,     --  input.wire
			output => bus_conversion6_output_wire  -- output.wire
		);

	ts_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => Ts,               --  input.wire
			output => ts_0_output_wire  -- output.wire
		);

	bus_conversion5 : component alt_dspbuilder_cast_GNLZYLEWIQ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast10_output_wire,          --  input.wire
			output => bus_conversion5_output_wire  -- output.wire
		);

	cast7 : component alt_dspbuilder_cast_GNSPENWJQH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vd_0_output_wire,  --  input.wire
			output => cast7_output_wire  -- output.wire
		);

	cast8 : component alt_dspbuilder_cast_GNQP67JAWW
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pll_3orden_change_pll_pi_z_1_sv2_0_e_wire, --  input.wire
			output => cast8_output_wire                          -- output.wire
		);

	cast9 : component alt_dspbuilder_cast_GNXY6JKR5E
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => wo_ref_0_output_wire, --  input.wire
			output => cast9_output_wire     -- output.wire
		);

	cast10 : component alt_dspbuilder_cast_GNRB4ECDTY
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pipelined_adder_result_wire, --  input.wire
			output => cast10_output_wire           -- output.wire
		);

	cast11 : component alt_dspbuilder_cast_GNCDTXOZMF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pipelined_adder1_result_wire, --  input.wire
			output => cast11_output_wire            -- output.wire
		);

	cast12 : component alt_dspbuilder_cast_GNWHGOINAS
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => x0_5_output_wire,   --  input.wire
			output => cast12_output_wire  -- output.wire
		);

end architecture rtl; -- of PLL_3orden_change_GN_PLL_3orden_change_PLL_PI_z
