-- PLL_3orden_change_GN.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PLL_3orden_change_GN is
	port (
		PLL_3orden_change_PLL_Vb_12b  : out std_logic_vector(11 downto 0);                    --  PLL_3orden_change_PLL_Vb_12b.wire
		clk60KPLL                     : in  std_logic                     := '0';             --                     clk60KPLL.wire
		Clock                         : in  std_logic                     := '0';             --                         Clock.clk
		aclr                          : in  std_logic                     := '0';             --                              .reset_n
		PLL_3orden_change_PLL_Va_12b  : out std_logic_vector(11 downto 0);                    --  PLL_3orden_change_PLL_Va_12b.wire
		PLL_3orden_change_PLL_Vm_12b  : out std_logic_vector(11 downto 0);                    --  PLL_3orden_change_PLL_Vm_12b.wire
		PLL_3orden_change_PLL_Vin_12b : out std_logic_vector(11 downto 0);                    -- PLL_3orden_change_PLL_Vin_12b.wire
		vin                           : in  std_logic_vector(11 downto 0) := (others => '0'); --                           vin.wire
		wot                           : out std_logic_vector(9 downto 0)                      --                           wot.wire
	);
end entity PLL_3orden_change_GN;

architecture rtl of PLL_3orden_change_GN is
	component alt_dspbuilder_clock_GNF343OQUJ is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNF343OQUJ;

	component PLL_3orden_change_GN_PLL_3orden_change_PLL is
		port (
			Vd      : out std_logic_vector(13 downto 0);                    -- wire
			Va_12b  : out std_logic_vector(11 downto 0);                    -- wire
			Vb_12b  : out std_logic_vector(11 downto 0);                    -- wire
			vit     : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wire
			Vin_12b : out std_logic_vector(11 downto 0);                    -- wire
			wot     : out std_logic_vector(9 downto 0);                     -- wire
			Vm_9b   : out std_logic_vector(8 downto 0);                     -- wire
			Clock   : in  std_logic                     := 'X';             -- clk
			aclr    : in  std_logic                     := 'X';             -- reset
			clk_60K : in  std_logic                     := 'X';             -- wire
			Vm_12b  : out std_logic_vector(11 downto 0)                     -- wire
		);
	end component PLL_3orden_change_GN_PLL_3orden_change_PLL;

	component alt_dspbuilder_port_GN4K6H3QBP is
		port (
			input  : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(11 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GN4K6H3QBP;

	component alt_dspbuilder_port_GNSSYS4J5R is
		port (
			input  : in  std_logic_vector(9 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(9 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNSSYS4J5R;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	signal clk60kpll_0_output_wire          : std_logic;                     -- clk60KPLL_0:output -> PLL_3orden_change_PLL_0:clk_60K
	signal vin_0_output_wire                : std_logic_vector(11 downto 0); -- vin_0:output -> PLL_3orden_change_PLL_0:vit
	signal pll_3orden_change_pll_0_wot_wire : std_logic_vector(9 downto 0);  -- PLL_3orden_change_PLL_0:wot -> wot_0:input
	signal clock_0_clock_output_clk         : std_logic;                     -- Clock_0:clock_out -> PLL_3orden_change_PLL_0:Clock
	signal clock_0_clock_output_reset       : std_logic;                     -- Clock_0:aclr_out -> PLL_3orden_change_PLL_0:aclr

begin

	clock_0 : component alt_dspbuilder_clock_GNF343OQUJ
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr_n    => aclr                        --             .reset_n
		);

	pll_3orden_change_pll_0 : component PLL_3orden_change_GN_PLL_3orden_change_PLL
		port map (
			Vd      => open,                             --      Vd.wire
			Va_12b  => PLL_3orden_change_PLL_Va_12b,     --  Va_12b.wire
			Vb_12b  => PLL_3orden_change_PLL_Vb_12b,     --  Vb_12b.wire
			vit     => vin_0_output_wire,                --     vit.wire
			Vin_12b => PLL_3orden_change_PLL_Vin_12b,    -- Vin_12b.wire
			wot     => pll_3orden_change_pll_0_wot_wire, --     wot.wire
			Vm_9b   => open,                             --   Vm_9b.wire
			Clock   => clock_0_clock_output_clk,         --   Clock.clk
			aclr    => clock_0_clock_output_reset,       --        .reset
			clk_60K => clk60kpll_0_output_wire,          -- clk_60K.wire
			Vm_12b  => PLL_3orden_change_PLL_Vm_12b      --  Vm_12b.wire
		);

	vin_0 : component alt_dspbuilder_port_GN4K6H3QBP
		port map (
			input  => vin,               --  input.wire
			output => vin_0_output_wire  -- output.wire
		);

	wot_0 : component alt_dspbuilder_port_GNSSYS4J5R
		port map (
			input  => pll_3orden_change_pll_0_wot_wire, --  input.wire
			output => wot                               -- output.wire
		);

	clk60kpll_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => clk60KPLL,               --  input.wire
			output => clk60kpll_0_output_wire  -- output.wire
		);

end architecture rtl; -- of PLL_3orden_change_GN
