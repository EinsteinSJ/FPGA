-- PLL_3orden_change_GN_PLL_3orden_change_PLL_IntegradorW_Comparador.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PLL_3orden_change_GN_PLL_3orden_change_PLL_IntegradorW_Comparador is
	port (
		Z     : out std_logic_vector(31 downto 0);                    --     Z.wire
		X     : in  std_logic_vector(31 downto 0) := (others => '0'); --     X.wire
		Y     : in  std_logic_vector(31 downto 0) := (others => '0'); --     Y.wire
		SAT   : out std_logic;                                        --   SAT.wire
		Clock : in  std_logic                     := '0';             -- Clock.clk
		aclr  : in  std_logic                     := '0'              --      .reset
	);
end entity PLL_3orden_change_GN_PLL_3orden_change_PLL_IntegradorW_Comparador;

architecture rtl of PLL_3orden_change_GN_PLL_3orden_change_PLL_IntegradorW_Comparador is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_multiplexer_GN2HWDO7FZ is
		generic (
			number_inputs          : natural  := 4;
			pipeline               : natural  := 0;
			width                  : positive := 8;
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(31 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(31 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GN2HWDO7FZ;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component alt_dspbuilder_pipelined_adder_GNY2JEH574 is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNY2JEH574;

	component alt_dspbuilder_comparator_GN is
		generic (
			Operator  : string  := "Altaeb";
			lpm_width : natural := 8
		);
		port (
			clock  : in  std_logic                              := 'X';             -- clk
			dataa  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			datab  : in  std_logic_vector(lpm_width-1 downto 0) := (others => 'X'); -- wire
			result : out std_logic;                                                 -- wire
			sclr   : in  std_logic                              := 'X'              -- clk
		);
	end component alt_dspbuilder_comparator_GN;

	component alt_dspbuilder_cast_GN46N4UJ5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic                    := 'X'; -- wire
			output : out std_logic_vector(0 downto 0)         -- wire
		);
	end component alt_dspbuilder_cast_GN46N4UJ5S;

	signal multiplexeruser_aclrgnd_output_wire      : std_logic;                     -- Multiplexeruser_aclrGND:output -> Multiplexer:user_aclr
	signal multiplexerenavcc_output_wire            : std_logic;                     -- MultiplexerenaVCC:output -> Multiplexer:ena
	signal pipelined_adder4user_aclrgnd_output_wire : std_logic;                     -- Pipelined_Adder4user_aclrGND:output -> Pipelined_Adder4:user_aclr
	signal pipelined_adder4enavcc_output_wire       : std_logic;                     -- Pipelined_Adder4enaVCC:output -> Pipelined_Adder4:ena
	signal x_0_output_wire                          : std_logic_vector(31 downto 0); -- X_0:output -> [Comparator:dataa, Multiplexer:in0, Pipelined_Adder4:dataa]
	signal y_0_output_wire                          : std_logic_vector(31 downto 0); -- Y_0:output -> [Comparator:datab, Pipelined_Adder4:datab]
	signal pipelined_adder4_result_wire             : std_logic_vector(31 downto 0); -- Pipelined_Adder4:result -> Multiplexer:in1
	signal multiplexer_result_wire                  : std_logic_vector(31 downto 0); -- Multiplexer:result -> Z_0:input
	signal comparator_result_wire                   : std_logic;                     -- Comparator:result -> [SAT_0:input, cast36:input]
	signal cast36_output_wire                       : std_logic_vector(0 downto 0);  -- cast36:output -> Multiplexer:sel
	signal clock_0_clock_output_clk                 : std_logic;                     -- Clock_0:clock_out -> [Comparator:clock, Multiplexer:clock, Pipelined_Adder4:clock]
	signal clock_0_clock_output_reset               : std_logic;                     -- Clock_0:aclr_out -> [Comparator:sclr, Multiplexer:aclr, Pipelined_Adder4:aclr]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	multiplexer : component alt_dspbuilder_multiplexer_GN2HWDO7FZ
		generic map (
			number_inputs          => 2,
			pipeline               => 0,
			width                  => 32,
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			sel       => cast36_output_wire,                  --        sel.wire
			result    => multiplexer_result_wire,             --     result.wire
			ena       => multiplexerenavcc_output_wire,       --        ena.wire
			user_aclr => multiplexeruser_aclrgnd_output_wire, --  user_aclr.wire
			in0       => x_0_output_wire,                     --        in0.wire
			in1       => pipelined_adder4_result_wire         --        in1.wire
		);

	multiplexeruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexeruser_aclrgnd_output_wire  -- output.wire
		);

	multiplexerenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexerenavcc_output_wire  -- output.wire
		);

	sat_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => comparator_result_wire, --  input.wire
			output => SAT                     -- output.wire
		);

	x_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => X,               --  input.wire
			output => x_0_output_wire  -- output.wire
		);

	pipelined_adder4 : component alt_dspbuilder_pipelined_adder_GNY2JEH574
		generic map (
			pipeline => 0,
			width    => 32
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => x_0_output_wire,                          --      dataa.wire
			datab     => y_0_output_wire,                          --      datab.wire
			result    => pipelined_adder4_result_wire,             --     result.wire
			user_aclr => pipelined_adder4user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder4enavcc_output_wire        --        ena.wire
		);

	pipelined_adder4user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder4user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder4enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder4enavcc_output_wire  -- output.wire
		);

	y_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => Y,               --  input.wire
			output => y_0_output_wire  -- output.wire
		);

	z_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => multiplexer_result_wire, --  input.wire
			output => Z                        -- output.wire
		);

	comparator : component alt_dspbuilder_comparator_GN
		generic map (
			Operator  => "Altageb",
			lpm_width => 32
		)
		port map (
			clock  => clock_0_clock_output_clk,   -- clock_sclr.clk
			sclr   => clock_0_clock_output_reset, --           .reset
			dataa  => x_0_output_wire,            --      dataa.wire
			datab  => y_0_output_wire,            --      datab.wire
			result => comparator_result_wire      --     result.wire
		);

	cast36 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => comparator_result_wire, --  input.wire
			output => cast36_output_wire      -- output.wire
		);

end architecture rtl; -- of PLL_3orden_change_GN_PLL_3orden_change_PLL_IntegradorW_Comparador
