-- PLL_3orden_change_GN_PLL_3orden_change_PLL_1erCon.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PLL_3orden_change_GN_PLL_3orden_change_PLL_1erCon is
	port (
		Clock      : in  std_logic                     := '0';             --      Clock.clk
		aclr       : in  std_logic                     := '0';             --           .reset
		id_14sfVin : out std_logic_vector(13 downto 0);                    -- id_14sfVin.wire
		Vin12b     : out std_logic_vector(11 downto 0);                    --     Vin12b.wire
		Vr         : in  std_logic_vector(11 downto 0) := (others => '0')  --         Vr.wire
	);
end entity PLL_3orden_change_GN_PLL_3orden_change_PLL_1erCon;

architecture rtl of PLL_3orden_change_GN_PLL_3orden_change_PLL_1erCon is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_cast_GNTSUCRN4Q is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNTSUCRN4Q;

	component alt_dspbuilder_cast_GNUYRTQ4QH is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNUYRTQ4QH;

	component alt_dspbuilder_cast_GNBZULANAF is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNBZULANAF;

	component alt_dspbuilder_cast_GNDS5WH6UV is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(11 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNDS5WH6UV;

	component alt_dspbuilder_constant_GNGPCXCFCV is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(12 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNGPCXCFCV;

	component alt_dspbuilder_pipelined_adder_GNY2JEH574 is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNY2JEH574;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_port_GNBOOX3JQY is
		port (
			input  : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNBOOX3JQY;

	component alt_dspbuilder_port_GN4K6H3QBP is
		port (
			input  : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(11 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GN4K6H3QBP;

	component alt_dspbuilder_cast_GNA5AA6QPF is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(12 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(12 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNA5AA6QPF;

	component alt_dspbuilder_cast_GN3AOOCYLL is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(11 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(12 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN3AOOCYLL;

	component alt_dspbuilder_cast_GN2UCHVFFC is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN2UCHVFFC;

	component alt_dspbuilder_cast_GN2YIIM3UI is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(12 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN2YIIM3UI;

	component alt_dspbuilder_cast_GNEX3PNEW7 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(12 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(11 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNEX3PNEW7;

	signal pipelined_adderuser_aclrgnd_output_wire : std_logic;                     -- Pipelined_Adderuser_aclrGND:output -> Pipelined_Adder:user_aclr
	signal pipelined_adderenavcc_output_wire       : std_logic;                     -- Pipelined_AdderenaVCC:output -> Pipelined_Adder:ena
	signal bus_conversion_output_wire              : std_logic_vector(23 downto 0); -- Bus_Conversion:output -> Binary_Point_Casting1:input
	signal binary_point_casting_output_wire        : std_logic_vector(12 downto 0); -- Binary_Point_Casting:output -> Pipelined_Adder:dataa
	signal cte_output_wire                         : std_logic_vector(12 downto 0); -- CTE:output -> Pipelined_Adder:datab
	signal bus_conversion3_output_wire             : std_logic_vector(13 downto 0); -- Bus_Conversion3:output -> id_14sfVin_0:input
	signal bus_conversion1_output_wire             : std_logic_vector(11 downto 0); -- Bus_Conversion1:output -> Vin12b_0:input
	signal vr_0_output_wire                        : std_logic_vector(11 downto 0); -- Vr_0:output -> cast31:input
	signal cast31_output_wire                      : std_logic_vector(12 downto 0); -- cast31:output -> Binary_Point_Casting:input
	signal binary_point_casting1_output_wire       : std_logic_vector(23 downto 0); -- Binary_Point_Casting1:output -> cast32:input
	signal cast32_output_wire                      : std_logic_vector(13 downto 0); -- cast32:output -> Bus_Conversion3:input
	signal pipelined_adder_result_wire             : std_logic_vector(12 downto 0); -- Pipelined_Adder:result -> [cast33:input, cast34:input]
	signal cast33_output_wire                      : std_logic_vector(23 downto 0); -- cast33:output -> Bus_Conversion:input
	signal cast34_output_wire                      : std_logic_vector(11 downto 0); -- cast34:output -> Bus_Conversion1:input
	signal clock_0_clock_output_clk                : std_logic;                     -- Clock_0:clock_out -> Pipelined_Adder:clock
	signal clock_0_clock_output_reset              : std_logic;                     -- Clock_0:aclr_out -> Pipelined_Adder:aclr

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	bus_conversion3 : component alt_dspbuilder_cast_GNTSUCRN4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast32_output_wire,          --  input.wire
			output => bus_conversion3_output_wire  -- output.wire
		);

	binary_point_casting1 : component alt_dspbuilder_cast_GNUYRTQ4QH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => bus_conversion_output_wire,        --  input.wire
			output => binary_point_casting1_output_wire  -- output.wire
		);

	bus_conversion : component alt_dspbuilder_cast_GNBZULANAF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast33_output_wire,         --  input.wire
			output => bus_conversion_output_wire  -- output.wire
		);

	bus_conversion1 : component alt_dspbuilder_cast_GNDS5WH6UV
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast34_output_wire,          --  input.wire
			output => bus_conversion1_output_wire  -- output.wire
		);

	cte : component alt_dspbuilder_constant_GNGPCXCFCV
		generic map (
			BitPattern => "0011101011111",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 13
		)
		port map (
			output => cte_output_wire  -- output.wire
		);

	pipelined_adder : component alt_dspbuilder_pipelined_adder_GNY2JEH574
		generic map (
			pipeline => 0,
			width    => 13
		)
		port map (
			clock     => clock_0_clock_output_clk,                -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,              --           .reset
			dataa     => binary_point_casting_output_wire,        --      dataa.wire
			datab     => cte_output_wire,                         --      datab.wire
			result    => pipelined_adder_result_wire,             --     result.wire
			user_aclr => pipelined_adderuser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adderenavcc_output_wire        --        ena.wire
		);

	pipelined_adderuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adderuser_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adderenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adderenavcc_output_wire  -- output.wire
		);

	id_14sfvin_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => bus_conversion3_output_wire, --  input.wire
			output => id_14sfVin                   -- output.wire
		);

	vr_0 : component alt_dspbuilder_port_GN4K6H3QBP
		port map (
			input  => Vr,               --  input.wire
			output => vr_0_output_wire  -- output.wire
		);

	vin12b_0 : component alt_dspbuilder_port_GN4K6H3QBP
		port map (
			input  => bus_conversion1_output_wire, --  input.wire
			output => Vin12b                       -- output.wire
		);

	binary_point_casting : component alt_dspbuilder_cast_GNA5AA6QPF
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast31_output_wire,               --  input.wire
			output => binary_point_casting_output_wire  -- output.wire
		);

	cast31 : component alt_dspbuilder_cast_GN3AOOCYLL
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vr_0_output_wire,   --  input.wire
			output => cast31_output_wire  -- output.wire
		);

	cast32 : component alt_dspbuilder_cast_GN2UCHVFFC
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => binary_point_casting1_output_wire, --  input.wire
			output => cast32_output_wire                 -- output.wire
		);

	cast33 : component alt_dspbuilder_cast_GN2YIIM3UI
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pipelined_adder_result_wire, --  input.wire
			output => cast33_output_wire           -- output.wire
		);

	cast34 : component alt_dspbuilder_cast_GNEX3PNEW7
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pipelined_adder_result_wire, --  input.wire
			output => cast34_output_wire           -- output.wire
		);

end architecture rtl; -- of PLL_3orden_change_GN_PLL_3orden_change_PLL_1erCon
