-- PLL_3orden_change_GN_PLL_3orden_change_PLL_SOGI.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PLL_3orden_change_GN_PLL_3orden_change_PLL_SOGI is
	port (
		Va      : out std_logic_vector(13 downto 0);                    --      Va.wire
		wo      : in  std_logic_vector(17 downto 0) := (others => '0'); --      wo.wire
		Vin     : in  std_logic_vector(13 downto 0) := (others => '0'); --     Vin.wire
		Vb      : out std_logic_vector(13 downto 0);                    --      Vb.wire
		Clk_60K : in  std_logic                     := '0';             -- Clk_60K.wire
		Clock   : in  std_logic                     := '0';             --   Clock.clk
		aclr    : in  std_logic                     := '0';             --        .reset
		Ts      : in  std_logic_vector(31 downto 0) := (others => '0')  --      Ts.wire
	);
end entity PLL_3orden_change_GN_PLL_3orden_change_PLL_SOGI;

architecture rtl of PLL_3orden_change_GN_PLL_3orden_change_PLL_SOGI is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_multiplier_GNER2DIGMG is
		generic (
			aWidth                         : natural := 8;
			Signed                         : natural := 0;
			bWidth                         : natural := 8;
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			pipeline                       : integer := 0;
			OutputLsb                      : integer := 0;
			OutputMsb                      : integer := 8
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GNER2DIGMG;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_cast_GNTSUCRN4Q is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNTSUCRN4Q;

	component alt_dspbuilder_cast_GNXTVWHWB4 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNXTVWHWB4;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_pipelined_adder_GNY2JEH574 is
		generic (
			pipeline : integer := 0;
			width    : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNY2JEH574;

	component alt_dspbuilder_port_GNBOOX3JQY is
		port (
			input  : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNBOOX3JQY;

	component alt_dspbuilder_port_GN2CABCRLL is
		port (
			input  : in  std_logic_vector(17 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(17 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GN2CABCRLL;

	component PLL_3orden_change_GN_PLL_3orden_change_PLL_SOGI_1_sv2 is
		port (
			CLK_60K : in  std_logic                     := 'X';             -- wire
			Out1    : out std_logic_vector(31 downto 0);                    -- wire
			In_1    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			Ts      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			Clock   : in  std_logic                     := 'X';             -- clk
			aclr    : in  std_logic                     := 'X'              -- reset
		);
	end component PLL_3orden_change_GN_PLL_3orden_change_PLL_SOGI_1_sv2;

	component PLL_3orden_change_GN_PLL_3orden_change_PLL_SOGI_1_sv1 is
		port (
			In_1    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			CLK_60K : in  std_logic                     := 'X';             -- wire
			Ts      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			Clock   : in  std_logic                     := 'X';             -- clk
			aclr    : in  std_logic                     := 'X';             -- reset
			Out1    : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component PLL_3orden_change_GN_PLL_3orden_change_PLL_SOGI_1_sv1;

	component alt_dspbuilder_cast_GNCWEIKWMJ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNCWEIKWMJ;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component alt_dspbuilder_cast_GNDI2FRQVQ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(17 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNDI2FRQVQ;

	signal multiplier1user_aclrgnd_output_wire          : std_logic;                     -- Multiplier1user_aclrGND:output -> Multiplier1:user_aclr
	signal multiplier1enavcc_output_wire                : std_logic;                     -- Multiplier1enaVCC:output -> Multiplier1:ena
	signal pipelined_adderuser_aclrgnd_output_wire      : std_logic;                     -- Pipelined_Adderuser_aclrGND:output -> Pipelined_Adder:user_aclr
	signal pipelined_adderenavcc_output_wire            : std_logic;                     -- Pipelined_AdderenaVCC:output -> Pipelined_Adder:ena
	signal multiplieruser_aclrgnd_output_wire           : std_logic;                     -- Multiplieruser_aclrGND:output -> Multiplier:user_aclr
	signal multiplierenavcc_output_wire                 : std_logic;                     -- MultiplierenaVCC:output -> Multiplier:ena
	signal pipelined_adder1user_aclrgnd_output_wire     : std_logic;                     -- Pipelined_Adder1user_aclrGND:output -> Pipelined_Adder1:user_aclr
	signal pipelined_adder1enavcc_output_wire           : std_logic;                     -- Pipelined_Adder1enaVCC:output -> Pipelined_Adder1:ena
	signal clk_60k_0_output_wire                        : std_logic;                     -- Clk_60K_0:output -> [PLL_3orden_change_PLL_SOGI_1_sv1_0:CLK_60K, PLL_3orden_change_PLL_SOGI_1_sv2_0:CLK_60K]
	signal ts_0_output_wire                             : std_logic_vector(31 downto 0); -- Ts_0:output -> [PLL_3orden_change_PLL_SOGI_1_sv1_0:Ts, PLL_3orden_change_PLL_SOGI_1_sv2_0:Ts]
	signal pll_3orden_change_pll_sogi_1_sv2_0_out1_wire : std_logic_vector(31 downto 0); -- PLL_3orden_change_PLL_SOGI_1_sv2_0:Out1 -> AltBus:input
	signal pll_3orden_change_pll_sogi_1_sv1_0_out1_wire : std_logic_vector(13 downto 0); -- PLL_3orden_change_PLL_SOGI_1_sv1_0:Out1 -> [AltBus1:input, Multiplier1:datab, Va_0:input]
	signal vin_0_output_wire                            : std_logic_vector(13 downto 0); -- Vin_0:output -> Bus_Conversion2:input
	signal bus_conversion6_output_wire                  : std_logic_vector(13 downto 0); -- Bus_Conversion6:output -> [Multiplier1:dataa, Multiplier:datab]
	signal multiplier_result_wire                       : std_logic_vector(15 downto 0); -- Multiplier:result -> PLL_3orden_change_PLL_SOGI_1_sv1_0:In_1
	signal multiplier1_result_wire                      : std_logic_vector(15 downto 0); -- Multiplier1:result -> PLL_3orden_change_PLL_SOGI_1_sv2_0:In_1
	signal bus_conversion2_output_wire                  : std_logic_vector(13 downto 0); -- Bus_Conversion2:output -> Pipelined_Adder:dataa
	signal altbus1_output_wire                          : std_logic_vector(13 downto 0); -- AltBus1:output -> Pipelined_Adder:datab
	signal pipelined_adder_result_wire                  : std_logic_vector(13 downto 0); -- Pipelined_Adder:result -> Pipelined_Adder1:dataa
	signal altbus_output_wire                           : std_logic_vector(13 downto 0); -- AltBus:output -> [Pipelined_Adder1:datab, Vb_0:input]
	signal pipelined_adder1_result_wire                 : std_logic_vector(13 downto 0); -- Pipelined_Adder1:result -> Multiplier:dataa
	signal wo_0_output_wire                             : std_logic_vector(17 downto 0); -- wo_0:output -> cast59:input
	signal cast59_output_wire                           : std_logic_vector(13 downto 0); -- cast59:output -> Bus_Conversion6:input
	signal clock_0_clock_output_clk                     : std_logic;                     -- Clock_0:clock_out -> [Multiplier1:clock, Multiplier:clock, PLL_3orden_change_PLL_SOGI_1_sv1_0:Clock, PLL_3orden_change_PLL_SOGI_1_sv2_0:Clock, Pipelined_Adder1:clock, Pipelined_Adder:clock]
	signal clock_0_clock_output_reset                   : std_logic;                     -- Clock_0:aclr_out -> [Multiplier1:aclr, Multiplier:aclr, PLL_3orden_change_PLL_SOGI_1_sv1_0:aclr, PLL_3orden_change_PLL_SOGI_1_sv2_0:aclr, Pipelined_Adder1:aclr, Pipelined_Adder:aclr]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	multiplier1 : component alt_dspbuilder_multiplier_GNER2DIGMG
		generic map (
			aWidth                         => 14,
			Signed                         => 1,
			bWidth                         => 14,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 1,
			OutputLsb                      => 10,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,                     -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,                   --           .reset
			dataa     => bus_conversion6_output_wire,                  --      dataa.wire
			datab     => pll_3orden_change_pll_sogi_1_sv1_0_out1_wire, --      datab.wire
			result    => multiplier1_result_wire,                      --     result.wire
			user_aclr => multiplier1user_aclrgnd_output_wire,          --  user_aclr.wire
			ena       => multiplier1enavcc_output_wire                 --        ena.wire
		);

	multiplier1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier1user_aclrgnd_output_wire  -- output.wire
		);

	multiplier1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplier1enavcc_output_wire  -- output.wire
		);

	bus_conversion2 : component alt_dspbuilder_cast_GNTSUCRN4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vin_0_output_wire,           --  input.wire
			output => bus_conversion2_output_wire  -- output.wire
		);

	altbus : component alt_dspbuilder_cast_GNXTVWHWB4
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pll_3orden_change_pll_sogi_1_sv2_0_out1_wire, --  input.wire
			output => altbus_output_wire                            -- output.wire
		);

	clk_60k_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => Clk_60K,               --  input.wire
			output => clk_60k_0_output_wire  -- output.wire
		);

	pipelined_adder : component alt_dspbuilder_pipelined_adder_GNY2JEH574
		generic map (
			pipeline => 0,
			width    => 14
		)
		port map (
			clock     => clock_0_clock_output_clk,                -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,              --           .reset
			dataa     => bus_conversion2_output_wire,             --      dataa.wire
			datab     => altbus1_output_wire,                     --      datab.wire
			result    => pipelined_adder_result_wire,             --     result.wire
			user_aclr => pipelined_adderuser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adderenavcc_output_wire        --        ena.wire
		);

	pipelined_adderuser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adderuser_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adderenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adderenavcc_output_wire  -- output.wire
		);

	va_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => pll_3orden_change_pll_sogi_1_sv1_0_out1_wire, --  input.wire
			output => Va                                            -- output.wire
		);

	vb_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => altbus_output_wire, --  input.wire
			output => Vb                  -- output.wire
		);

	wo_0 : component alt_dspbuilder_port_GN2CABCRLL
		port map (
			input  => wo,               --  input.wire
			output => wo_0_output_wire  -- output.wire
		);

	altbus1 : component alt_dspbuilder_cast_GNTSUCRN4Q
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pll_3orden_change_pll_sogi_1_sv1_0_out1_wire, --  input.wire
			output => altbus1_output_wire                           -- output.wire
		);

	multiplier : component alt_dspbuilder_multiplier_GNER2DIGMG
		generic map (
			aWidth                         => 14,
			Signed                         => 1,
			bWidth                         => 14,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 1,
			OutputLsb                      => 10,
			OutputMsb                      => 25
		)
		port map (
			clock     => clock_0_clock_output_clk,           -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,         --           .reset
			dataa     => pipelined_adder1_result_wire,       --      dataa.wire
			datab     => bus_conversion6_output_wire,        --      datab.wire
			result    => multiplier_result_wire,             --     result.wire
			user_aclr => multiplieruser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => multiplierenavcc_output_wire        --        ena.wire
		);

	multiplieruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplieruser_aclrgnd_output_wire  -- output.wire
		);

	multiplierenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplierenavcc_output_wire  -- output.wire
		);

	vin_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => Vin,               --  input.wire
			output => vin_0_output_wire  -- output.wire
		);

	pll_3orden_change_pll_sogi_1_sv2_0 : component PLL_3orden_change_GN_PLL_3orden_change_PLL_SOGI_1_sv2
		port map (
			CLK_60K => clk_60k_0_output_wire,                        -- CLK_60K.wire
			Out1    => pll_3orden_change_pll_sogi_1_sv2_0_out1_wire, --    Out1.wire
			In_1    => multiplier1_result_wire,                      --    In_1.wire
			Ts      => ts_0_output_wire,                             --      Ts.wire
			Clock   => clock_0_clock_output_clk,                     --   Clock.clk
			aclr    => clock_0_clock_output_reset                    --        .reset
		);

	pll_3orden_change_pll_sogi_1_sv1_0 : component PLL_3orden_change_GN_PLL_3orden_change_PLL_SOGI_1_sv1
		port map (
			In_1    => multiplier_result_wire,                       --    In_1.wire
			CLK_60K => clk_60k_0_output_wire,                        -- CLK_60K.wire
			Ts      => ts_0_output_wire,                             --      Ts.wire
			Clock   => clock_0_clock_output_clk,                     --   Clock.clk
			aclr    => clock_0_clock_output_reset,                   --        .reset
			Out1    => pll_3orden_change_pll_sogi_1_sv1_0_out1_wire  --    Out1.wire
		);

	pipelined_adder1 : component alt_dspbuilder_pipelined_adder_GNY2JEH574
		generic map (
			pipeline => 0,
			width    => 14
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => pipelined_adder_result_wire,              --      dataa.wire
			datab     => altbus_output_wire,                       --      datab.wire
			result    => pipelined_adder1_result_wire,             --     result.wire
			user_aclr => pipelined_adder1user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder1enavcc_output_wire        --        ena.wire
		);

	pipelined_adder1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder1user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder1enavcc_output_wire  -- output.wire
		);

	bus_conversion6 : component alt_dspbuilder_cast_GNCWEIKWMJ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast59_output_wire,          --  input.wire
			output => bus_conversion6_output_wire  -- output.wire
		);

	ts_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => Ts,               --  input.wire
			output => ts_0_output_wire  -- output.wire
		);

	cast59 : component alt_dspbuilder_cast_GNDI2FRQVQ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => wo_0_output_wire,   --  input.wire
			output => cast59_output_wire  -- output.wire
		);

end architecture rtl; -- of PLL_3orden_change_GN_PLL_3orden_change_PLL_SOGI
