-- PLL_3orden_change_GN_PLL_3orden_change_PLL_Vm_Num.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PLL_3orden_change_GN_PLL_3orden_change_PLL_Vm_Num is
	port (
		Vmi   : in  std_logic_vector(14 downto 0) := (others => '0'); --   Vmi.wire
		Clock : in  std_logic                     := '0';             -- Clock.clk
		aclr  : in  std_logic                     := '0';             --      .reset
		Vmo   : out std_logic_vector(8 downto 0)                      --   Vmo.wire
	);
end entity PLL_3orden_change_GN_PLL_3orden_change_PLL_Vm_Num;

architecture rtl of PLL_3orden_change_GN_PLL_3orden_change_PLL_Vm_Num is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_constant_GNQ42UAUVX is
		generic (
			BitPattern : string  := "0000";
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(12 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNQ42UAUVX;

	component alt_dspbuilder_port_GNIF77H5YS is
		port (
			input  : in  std_logic_vector(14 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(14 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNIF77H5YS;

	component alt_dspbuilder_multiplier_GNM7I5EZ6T is
		generic (
			aWidth                         : natural := 8;
			Signed                         : natural := 0;
			bWidth                         : natural := 8;
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			pipeline                       : integer := 0;
			OutputLsb                      : integer := 0;
			OutputMsb                      : integer := 8
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GNM7I5EZ6T;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_round_GNQI7H3AHU is
		generic (
			OUT_WIDTH_g     : natural := 6;
			IN_WIDTH_g      : natural := 8;
			PIPELINE_g      : natural := 0;
			ROUNDING_TYPE_g : string  := "TRUNCATE_LOW";
			SIGNED_g        : natural := 1
		);
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- wire
			datain    : in  std_logic_vector(10 downto 0) := (others => 'X'); -- wire
			dataout   : out std_logic_vector(8 downto 0);                     -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X'              -- wire
		);
	end component alt_dspbuilder_round_GNQI7H3AHU;

	component alt_dspbuilder_port_GNJVFJM3AT is
		port (
			input  : in  std_logic_vector(8 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(8 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNJVFJM3AT;

	component alt_dspbuilder_cast_GNN7MLWJTA is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(14 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNN7MLWJTA;

	signal multiplieruser_aclrgnd_output_wire : std_logic;                     -- Multiplieruser_aclrGND:output -> Multiplier:user_aclr
	signal multiplierenavcc_output_wire       : std_logic;                     -- MultiplierenaVCC:output -> Multiplier:ena
	signal rounduser_aclrgnd_output_wire      : std_logic;                     -- Rounduser_aclrGND:output -> Round:user_aclr
	signal roundresetgnd_output_wire          : std_logic;                     -- RoundresetGND:output -> Round:reset
	signal roundenavcc_output_wire            : std_logic;                     -- RoundenaVCC:output -> Round:ena
	signal multiplier_result_wire             : std_logic_vector(10 downto 0); -- Multiplier:result -> Round:datain
	signal sca_output_wire                    : std_logic_vector(12 downto 0); -- SCA:output -> Multiplier:datab
	signal round_dataout_wire                 : std_logic_vector(8 downto 0);  -- Round:dataout -> Vmo_0:input
	signal vmi_0_output_wire                  : std_logic_vector(14 downto 0); -- Vmi_0:output -> cast35:input
	signal cast35_output_wire                 : std_logic_vector(13 downto 0); -- cast35:output -> Multiplier:dataa
	signal clock_0_clock_output_clk           : std_logic;                     -- Clock_0:clock_out -> [Multiplier:clock, Round:clk]
	signal clock_0_clock_output_reset         : std_logic;                     -- Clock_0:aclr_out -> [Multiplier:aclr, Round:reset]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	sca : component alt_dspbuilder_constant_GNQ42UAUVX
		generic map (
			BitPattern => "1110100101011",
			HDLTYPE    => "STD_LOGIC_VECTOR",
			width      => 13
		)
		port map (
			output => sca_output_wire  -- output.wire
		);

	vmi_0 : component alt_dspbuilder_port_GNIF77H5YS
		port map (
			input  => Vmi,               --  input.wire
			output => vmi_0_output_wire  -- output.wire
		);

	multiplier : component alt_dspbuilder_multiplier_GNM7I5EZ6T
		generic map (
			aWidth                         => 14,
			Signed                         => 0,
			bWidth                         => 13,
			DEDICATED_MULTIPLIER_CIRCUITRY => "NO",
			pipeline                       => 1,
			OutputLsb                      => 14,
			OutputMsb                      => 24
		)
		port map (
			clock     => clock_0_clock_output_clk,           -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,         --           .reset
			dataa     => cast35_output_wire,                 --      dataa.wire
			datab     => sca_output_wire,                    --      datab.wire
			result    => multiplier_result_wire,             --     result.wire
			user_aclr => multiplieruser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => multiplierenavcc_output_wire        --        ena.wire
		);

	multiplieruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplieruser_aclrgnd_output_wire  -- output.wire
		);

	multiplierenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplierenavcc_output_wire  -- output.wire
		);

	round : component alt_dspbuilder_round_GNQI7H3AHU
		generic map (
			OUT_WIDTH_g     => 9,
			IN_WIDTH_g      => 11,
			PIPELINE_g      => 0,
			ROUNDING_TYPE_g => "TRUNCATE_LOW",
			SIGNED_g        => 0
		)
		port map (
			clk       => clock_0_clock_output_clk,      -- clk_reset.clk
			reset     => clock_0_clock_output_reset,    --          .reset
			datain    => multiplier_result_wire,        --    datain.wire
			dataout   => round_dataout_wire,            --   dataout.wire
			ena       => roundenavcc_output_wire,       --       ena.wire
			user_aclr => rounduser_aclrgnd_output_wire  -- user_aclr.wire
		);

	rounduser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => rounduser_aclrgnd_output_wire  -- output.wire
		);

	roundresetgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => roundresetgnd_output_wire  -- output.wire
		);

	roundenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => roundenavcc_output_wire  -- output.wire
		);

	vmo_0 : component alt_dspbuilder_port_GNJVFJM3AT
		port map (
			input  => round_dataout_wire, --  input.wire
			output => Vmo                 -- output.wire
		);

	cast35 : component alt_dspbuilder_cast_GNN7MLWJTA
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vmi_0_output_wire,  --  input.wire
			output => cast35_output_wire  -- output.wire
		);

end architecture rtl; -- of PLL_3orden_change_GN_PLL_3orden_change_PLL_Vm_Num
