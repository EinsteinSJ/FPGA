-- PLL_3orden_change_GN_PLL_3orden_change_PLL_Signals.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity PLL_3orden_change_GN_PLL_3orden_change_PLL_Signals is
	port (
		Clock : in  std_logic                     := '0';             -- Clock.clk
		aclr  : in  std_logic                     := '0';             --      .reset
		Vm    : in  std_logic_vector(14 downto 0) := (others => '0'); --    Vm.wire
		Vb    : in  std_logic_vector(13 downto 0) := (others => '0'); --    Vb.wire
		Vin   : in  std_logic_vector(13 downto 0) := (others => '0'); --   Vin.wire
		Vb_2  : out std_logic_vector(21 downto 0);                    --  Vb_2.wire
		Vin_2 : out std_logic_vector(21 downto 0);                    -- Vin_2.wire
		Va_2  : out std_logic_vector(21 downto 0);                    --  Va_2.wire
		Va    : in  std_logic_vector(13 downto 0) := (others => '0'); --    Va.wire
		Vm_2  : out std_logic_vector(21 downto 0)                     --  Vm_2.wire
	);
end entity PLL_3orden_change_GN_PLL_3orden_change_PLL_Signals;

architecture rtl of PLL_3orden_change_GN_PLL_3orden_change_PLL_Signals is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_cast_GNNPYFJRPJ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(21 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(21 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNNPYFJRPJ;

	component alt_dspbuilder_port_GNBVD2CPQ4 is
		port (
			input  : in  std_logic_vector(21 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(21 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNBVD2CPQ4;

	component alt_dspbuilder_port_GNIF77H5YS is
		port (
			input  : in  std_logic_vector(14 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(14 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNIF77H5YS;

	component alt_dspbuilder_port_GNBOOX3JQY is
		port (
			input  : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(13 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNBOOX3JQY;

	component alt_dspbuilder_cast_GNMFPTKSML is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(13 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(21 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNMFPTKSML;

	component alt_dspbuilder_cast_GNM5FFDTMH is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(14 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(21 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNM5FFDTMH;

	signal bus_conversion_vin_output_wire : std_logic_vector(21 downto 0); -- Bus_Conversion_Vin:output -> Vin_2_0:input
	signal bus_conversion_va_output_wire  : std_logic_vector(21 downto 0); -- Bus_Conversion_Va:output -> Va_2_0:input
	signal bus_conversion_vb_output_wire  : std_logic_vector(21 downto 0); -- Bus_Conversion_Vb:output -> Vb_2_0:input
	signal bus_conversion_vb1_output_wire : std_logic_vector(21 downto 0); -- Bus_Conversion_Vb1:output -> Vm_2_0:input
	signal va_0_output_wire               : std_logic_vector(13 downto 0); -- Va_0:output -> cast15:input
	signal cast15_output_wire             : std_logic_vector(21 downto 0); -- cast15:output -> Bus_Conversion_Va:input
	signal vb_0_output_wire               : std_logic_vector(13 downto 0); -- Vb_0:output -> cast16:input
	signal cast16_output_wire             : std_logic_vector(21 downto 0); -- cast16:output -> Bus_Conversion_Vb:input
	signal vm_0_output_wire               : std_logic_vector(14 downto 0); -- Vm_0:output -> cast17:input
	signal cast17_output_wire             : std_logic_vector(21 downto 0); -- cast17:output -> Bus_Conversion_Vb1:input
	signal vin_0_output_wire              : std_logic_vector(13 downto 0); -- Vin_0:output -> cast18:input
	signal cast18_output_wire             : std_logic_vector(21 downto 0); -- cast18:output -> Bus_Conversion_Vin:input

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => open,  -- clock_output.clk
			aclr_out  => open,  --             .reset
			clock     => Clock, --        clock.clk
			aclr      => aclr   --             .reset
		);

	bus_conversion_vb1 : component alt_dspbuilder_cast_GNNPYFJRPJ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast17_output_wire,             --  input.wire
			output => bus_conversion_vb1_output_wire  -- output.wire
		);

	vm_2_0 : component alt_dspbuilder_port_GNBVD2CPQ4
		port map (
			input  => bus_conversion_vb1_output_wire, --  input.wire
			output => Vm_2                            -- output.wire
		);

	vin_2_0 : component alt_dspbuilder_port_GNBVD2CPQ4
		port map (
			input  => bus_conversion_vin_output_wire, --  input.wire
			output => Vin_2                           -- output.wire
		);

	bus_conversion_vb : component alt_dspbuilder_cast_GNNPYFJRPJ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast16_output_wire,            --  input.wire
			output => bus_conversion_vb_output_wire  -- output.wire
		);

	bus_conversion_va : component alt_dspbuilder_cast_GNNPYFJRPJ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast15_output_wire,            --  input.wire
			output => bus_conversion_va_output_wire  -- output.wire
		);

	va_2_0 : component alt_dspbuilder_port_GNBVD2CPQ4
		port map (
			input  => bus_conversion_va_output_wire, --  input.wire
			output => Va_2                           -- output.wire
		);

	vm_0 : component alt_dspbuilder_port_GNIF77H5YS
		port map (
			input  => Vm,               --  input.wire
			output => vm_0_output_wire  -- output.wire
		);

	vb_2_0 : component alt_dspbuilder_port_GNBVD2CPQ4
		port map (
			input  => bus_conversion_vb_output_wire, --  input.wire
			output => Vb_2                           -- output.wire
		);

	bus_conversion_vin : component alt_dspbuilder_cast_GNNPYFJRPJ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast18_output_wire,             --  input.wire
			output => bus_conversion_vin_output_wire  -- output.wire
		);

	vin_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => Vin,               --  input.wire
			output => vin_0_output_wire  -- output.wire
		);

	va_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => Va,               --  input.wire
			output => va_0_output_wire  -- output.wire
		);

	vb_0 : component alt_dspbuilder_port_GNBOOX3JQY
		port map (
			input  => Vb,               --  input.wire
			output => vb_0_output_wire  -- output.wire
		);

	cast15 : component alt_dspbuilder_cast_GNMFPTKSML
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => va_0_output_wire,   --  input.wire
			output => cast15_output_wire  -- output.wire
		);

	cast16 : component alt_dspbuilder_cast_GNMFPTKSML
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vb_0_output_wire,   --  input.wire
			output => cast16_output_wire  -- output.wire
		);

	cast17 : component alt_dspbuilder_cast_GNM5FFDTMH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vm_0_output_wire,   --  input.wire
			output => cast17_output_wire  -- output.wire
		);

	cast18 : component alt_dspbuilder_cast_GNMFPTKSML
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => vin_0_output_wire,  --  input.wire
			output => cast18_output_wire  -- output.wire
		);

end architecture rtl; -- of PLL_3orden_change_GN_PLL_3orden_change_PLL_Signals
